`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: X-Force Red
// Engineer: Grzegorz Wypych (h0rac)
// 
// Create Date: 10/21/2019 01:53:37 AM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module top(
  input clk_27,
  input rst_n,
  input ftdi_rx,
  input trigger_in,
  input gpio_in1,
  input gpio_in2,
  output gpio_out,
  output ftdi_tx,
  output led0_g,
  output led0_r,
  output led0_b,
  output led2_g,
  output led2_r,
  output led2_b,
  output led_blink,
  output led5_debug,
  output led6_debug,
  output debug_io0_14_p30,
  output led_glitch_out,
  output wire glitch_out,
  output invert_glitch_out,
  output wire reset_out
    );
 
//  assign target_tx = ftdi_rx;
//  assign target_rx = ftdi_tx;

parameter AUTO = 2'd2;

wire clk;
wire rst;

wire bit_out;
wire active;

wire [31:0] glitch_delay;
wire [31:0] glitch_width;
wire [31:0] glitch_count;
wire [31:0] glitch_gap;
wire [31:0] glitch_max;
wire [31:0] reset_target;
wire armed;
wire glitched;
wire finished;
wire vstart; // glitch_out startup value
wire invert_trigger;
wire [1:0] force_state;
wire reset_glitcher;

// counter for main loop
reg [31:0] counter;

pll100MHz PLL1(
  .clkout(), //output clkout
  .clkin(clk_27), //input clkin
  .clkoutd(clk)
);
assign rst = ~rst_n;

cmd cmd_inst
(
  .clk(clk),
  .rst(rst),
  .din(ftdi_rx),
  .dout(bit_out),
  .trigger_in(trigger_in),
  .glitch_delay(glitch_delay),
  .glitch_width(glitch_width),
  .glitch_count(glitch_count),
  .glitch_gap(glitch_gap),
  .glitch_max(glitch_max),
  .armed(armed),
  .finished(finished),
  .glitched(glitched),
  .glitch_out(glitch_out),
  .force_state(force_state),
  .reset_glitcher(reset_glitcher),
  .vstart(vstart),
  .invert_trigger(invert_trigger),
  .reset_target(reset_target),
  .gpio_in1(gpio_in1),
  .gpio_in2(gpio_in2),
  .gpio_out(gpio_out)
  );   
  assign ftdi_tx =  bit_out;
  assign gpio_out = gpio_out;
 
 // reset target feature
// assign rst_out = reset_target ? 1'b0 : 1'b1;
wire glitch;
wire trigger;
assign trigger = invert_trigger ^ trigger_in;
assign glitch_out = force_state != AUTO ? force_state : glitch;
assign invert_glitch_out = !glitch_out;
wire enable =  (force_state == AUTO && (((armed && !finished) && trigger) || (glitch_max && glitched && !finished)));
 
 glitch glitchi
 (
  .clk(clk),
  .rst(rst || reset_glitcher),
  .enable(enable),
  .vout(glitch),
  .glitch_delay(glitch_delay),
  .glitch_width(glitch_width),
  .glitch_count(glitch_count),
  .glitch_gap(glitch_gap),
  .glitch_max(glitch_max),
  .glitched(glitched),
  .vstart(vstart),
  .finished(finished),
  .reset_target(reset_target),
  .reset_out(reset_out)
 );
 
  // LD0 - BLUE armed, GREEN glitching started, RED finished
  
   pwm pwm_led0_r (
    .clk(clk),
    .duty(8'd64),
    .signal(finished),
    .state(led0_r)
   );
   
   pwm pwm_led0_g (
    .clk(clk),
    .duty(8'd16),
    .signal(glitched && !finished),
    .state(led0_g)
   );
   
   pwm pwm_led0_b (
    .clk(clk),
    .duty(8'd64),
    .signal(!glitched && armed),
    .state(led0_b)
   );

   // LD1 - 
   
//   pwm pwm_led1_r (
//    .clk(clk),
//    .duty(64),
//    .signal(armed),
//    .state(led1_r)
//   );
   
//   pwm pwm_led1_g (
//    .clk(clk),
//    .duty(64),
//    .signal(armed),
//    .state(led1_g)
//   );
             
//   pwm pwm_led1_b (
//    .clk(clk),
//    .duty(0),
//    .signal(0),
//    .state(led1_b)
//   );
   
   // LD2 - trigger
          
   pwm pwm_led2_r (
    .clk(clk),
    .duty(8'd32),
    .signal(trigger_in),
    .state(led2_r)
   );
   
   pwm pwm_led2_g (
    .clk(clk),
    .duty(8'd4),
    .signal(trigger_in),
    .state(led2_g)
   );
                      
   pwm pwm_led2_b (
    .clk(clk),
    .duty(8'd48),
    .signal(trigger_in),
    .state(led2_b)
   );

  //assign debug_enable = (armed && trigger_in) || (armed && !trigger_in_pullup);
  assign debug_io0_14_p30 = glitch_out;
  assign led5_debug = reset_out;
  assign led6_debug = reset_target;
  assign led_blink = counter[26];
  assign led_glitch_out = glitch_out;
  
  always @(posedge clk)
  begin
    counter <= counter + 1;
  end
 
endmodule
